module eight_bit_prio_enco(d_out, d_in);
   
   output [2:0] d_out;
   input [7:0] d_in;

   assign d_out = (d_in[0] ==1'b1) ? 3'b000:
                (d_in[1] ==1'b1) ? 3'b001:
                (d_in[2] ==1'b1) ? 3'b010:
                (d_in[3] ==1'b1) ? 3'b011:
                (d_in[4] ==1'b1) ? 3'b100:
                (d_in[5] ==1'b1 ) ? 3'b101:
                (d_in[6] ==1'b1 ) ? 3'b110:
                (d_in[7] ==1'b1 ) ? 3'b111 : 3'bxxx;

endmodule