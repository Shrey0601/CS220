`include "A2Q1_helper.v"
`include "A2Q1_gen_prop.v"
module eight_bit_lookahead_carry (
    carry_bus,cin,p,g
);
    output[8:1] carry_bus;
    input cin;
    input[8:1] p,g;
    helper h1(carry_bus[1],)
    for()
endmodule