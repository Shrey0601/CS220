module sequence_gen (
    in,clk,inputs
);
    output reg in;
    input clk;
    input 
endmodule